module and_g(input a,b,output y);

	y = assign(a&b);

endmodule
